`timescale 1ns / 1ps

import defines::*;

module tb_alu_control_unit;

endmodule
